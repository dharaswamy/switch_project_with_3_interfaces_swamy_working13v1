interface out_intf(input clk,rst);

logic read_0=1;
logic read_1=1;
logic read_2=1;
logic read_3=1;

logic ready_0;
logic ready_1;
logic ready_2;
logic  ready_3;

logic  [7:0] port_0;
logic  [7:0] port_1;
logic  [7:0] port_2;
logic [7:0] port_3;



endinterface:out_intf